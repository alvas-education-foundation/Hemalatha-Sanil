// Code your design here
module inverter (a, y);
  input a;
  output y;
  assign y=~a;
endmodule